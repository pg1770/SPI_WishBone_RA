`timescale 1ns / 1ps

module SPI_MASTER(
  input clk,
  input rst,
  output reg [40:0] data_out,
  input [40:0] data_in,
  output reg ack_out,
  input ack_in,
  output min,
  input mout
    );


endmodule
