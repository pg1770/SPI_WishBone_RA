`timescale 1ns / 1ps

module SPI_MASTER(
  input clk,
  input rst,
  output [40:0] bin,
  input [40:0] bout,
  output backin,
  input backout,
  output min,
  input mout
    );


endmodule
